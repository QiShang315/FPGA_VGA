`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/02/09 16:45:58
// Design Name: 
// Module Name: VGA_TOP
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

// TOP connects the Frame_Buffer and VGA_Sig_Gen modules, managing data flow and timing.
module VGA_TOP (
    input wire        CLK_100MHz,          // 100MHz clock input
    input wire        RESET,               // Reset signal

    // External data writing interface (e.g. CPU or external controller)
    //input wire [14:0] addr_A,             // д���ַ
    //input wire        data_in_A,          // д������ (1-bit)

    // VGA output signals
    output wire       VGA_HS,             // Horizontal sync signal
    output wire       VGA_VS,             // Vertical sync signal
    
    output wire [2:0] VGA_RED,           // Red colour output (3-bit)
    output wire [2:0] VGA_GREEN,        // Green colour output (3-bit)
    output wire [1:0] VGA_BLUE          // Blue colour output (2-bit)
);


   // Colour parameters: RED and BLUE definitions
   parameter RED_COLOR  = 16'hE003; // Definition for red colour
   parameter BLUE_COLOR = 16'h03E0; // Definition for blue colour


   wire DPR_CLK;   //25MHz clock from VGA_Sig_Gen

 // === 1Hz timer (25MHz / 25,000,000 = 1Hz) ===
    reg [24:0] sec_counter = 0;   // 25bit counter required (Max 33,554,432 > 25000000)
    reg toggle = 0;               // Toggle signal for swapping foreground and background colours


       always @(posedge DPR_CLK) begin
           if (RESET) begin
              sec_counter <= 0;
              toggle <= 0;
           end else if (sec_counter >= 25_000_000) begin  //Every time sec_counter reaches 25,000,000
             sec_counter <= 0;                           //Reset sec_counter to 0
             toggle <= ~toggle;                         //Flip the toggle signal (0 to 1 or 1 to 0) at 1Hz
          end else begin
             sec_counter <= sec_counter + 1;
           end
       end


   // Swap foreground and background colours
    wire [15:0] CONFIG_COLOURS;
    assign CONFIG_COLOURS = (toggle) ? RED_COLOR : BLUE_COLOR;  
  // If toggle is 1, use RED_COLOR for foreground,  BLUE_COLOR for background
  // If toggle is 0, use BLUE_COLOR for foreground,  RED_COLOR for background
       

 // Connect the Frame_Buffer and VGA_Sig_Gen modules
    wire [14:0] VGA_ADDR;    // Frame buffer address generated by VGA_Sig_Gen
    wire VGA_DATA;           // 1-bit pixel data read from the frame buffer for VGA

 // Port A (for data write operations)
    wire clk_A = CLK_100MHz;

 // Port B (for VGA read operations)
    wire clk_B = DPR_CLK;            // Read clock is the 25MHz clock provided by VGA_Sig_Gen
    wire [14:0] addr_B = VGA_ADDR;  // VGA read address generated by VGA_Sig_Gen
    wire data_out_B;               //  Frame_Buffe outout to VGA_Sig_Gen

// Instantiate the Frame_Buffer module (stores pixel data)
    Frame_Buffer frame_buffer_inst (
        .clk_A(clk_A),
        .addr_A(),
        .data_in_A(),
        .we_A(),
        .data_out_A(),  
        .clk_B(clk_B),          // DPR_CLK
        .addr_B(addr_B),        // VGA_ADDR
        .data_out_B(VGA_DATA)  // VGA_DATA
    );

// Instantiate the VGA_Sig_Gen module (generates VGA signals)
    VGA_Sig_Gen vga_sig_gen_inst (
        .CLK(CLK_100MHz),  
        .RESET(RESET),
        .CONFIG_COLOURS(CONFIG_COLOURS), 
        .DPR_CLK(DPR_CLK),
        .VGA_ADDR(VGA_ADDR),
        .VGA_DATA(VGA_DATA),
        .VGA_HS(VGA_HS),
        .VGA_VS(VGA_VS),
        .VGA_COLOUR({VGA_RED, VGA_GREEN, VGA_BLUE})
    );

endmodule